`ifndef __HAZARD_CONTROL_V__
`define __HAZARD_CONTROL_V__

`timescale 1ns/100ps

module hazard_detection (
    input is_branch,

    output if_flush,
    output id_flush,
);


endmodule

`endif // __HAZARD_CONTROL_V__